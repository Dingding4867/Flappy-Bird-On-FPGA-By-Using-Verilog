module DE1_SoC (CLOCK_50, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, KEY, LEDR, SW, GPIO_1);
	input logic CLOCK_50; // 50MHz clock.
	output logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
	output logic [9:0] LEDR;
	output logic [35:0] GPIO_1;
	input logic [3:0] KEY; // True when not pressed, False when pressed
	input logic [9:0] SW;
	
	logic reset;
	logic result;
	logic [31:0] div_clk;
	assign reset = SW[9];

	 
	 
	clock_divider cdiv (.clock(CLOCK_50),
							  .reset(reset),
							  .divided_clocks(div_clk));
							  
// Clock selection; allows for easy switching between simulation and board
// clocks
	logic clkSelect;
	// Uncomment ONE of the following two lines depending on intention
	
	
	//assign clkSelect = CLOCK_50; // for simulation
	assign clkSelect = div_clk[23]; // for pipe
	assign birdSelect = div_clk[14]; //  for bird
	assign userSelect = div_clk[14];
	assign computerSelect = div_clk[14];// for computer
	
	
		 /* Set up system base clock to 1526 Hz (50 MHz / 2**(14+1))
	    ===========================================================*/
	 logic [31:0] clk;
	 logic SYSTEM_CLOCK;
	 logic RST;
	 
	 clock_divider divider (.clock(CLOCK_50), .divided_clocks(clk));
	 
	 assign SYSTEM_CLOCK = clk[14]; // 1526 Hz clock signal	 
	 
	 assign RST = ~KEY[0];
	
	 
		 
	logic [15:0][15:0]RedPixels; // 16 x 16 array representing red LEDs
   logic [15:0][15:0]GrnPixels; // 16 x 16 array representing green LEDs 
	logic [3:0] fakeRandomPatterns;// 4-bit random number 16 possibilities, fake randoms
	logic [15:0] randomWall;// A single column(pipe) made up by random redPixels
	logic pressInput;
	logic death;// if the bird(Green) colide with the pipes(Red)
	logic [3:0] hundreds, tens, units;// 9-9-9 counters
	logic [6:0] HEX_0, HEX_1, HEX_2;
	logic constantDown;// bird constant down 1 pixel
	logic stablePressed;
	logic outofbounddeath;
	
	
	/* Standard LED Driver instantiation - set once and 'forget it'. 
	    See LEDDriver.sv for more info. Do not modify unless you know what you are doing! */
	LEDDriver Driver (.CLK(SYSTEM_CLOCK), .RST, .EnableCount(1'b1), .RedPixels, .GrnPixels, .GPIO_1);
	
	// These modules are dealing with pipes and their movement
	LFSR lfsr1 (.Clock(clkSelect), .Reset(reset), .patterns(fakeRandomPatterns));// generate the random number
	singleRandomColumn singleColumn (.Clock(clkSelect), .Reset(reset), .fakeRandom(fakeRandomPatterns), .wall(randomWall));// generate random clumn based on the random number generated by LFSR
	allPipes allColumn (.Clock(clkSelect), .Reset(reset | death | outofbounddeath), .randomPipes(randomWall), .RedPixels);// Control all pipes
	
	// These modules are dealing with bird(human controled)
	Userinput userinput (.Clock(userSelect), .Reset(reset), .key(~KEY[3]), .pressedKey(pressInput));
	Metastability meta (.in(pressInput), .Clock(userSelect), .out(stablePressed));
	Computerinput computerinput (.Clock(computerSelect), .Reset(reset), .tick(constantDown));
	
	edgeLight bound (.Clock(birdSelect), .Reset(reset| death| outofbounddeath),.upLight(GrnPixels[0][13]), .downLight(GrnPixels[15][13]), .up(stablePressed), .bottom(constantDown), .outDeath(outofbounddeath));
	
	normalLight normal0 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(1'b0), .nBottom(GrnPixels[1][13]), .lightOn(GrnPixels[0][13]));//0
	normalLight normal1 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[0][13]), .nBottom(GrnPixels[2][13]), .lightOn(GrnPixels[1][13]));
	normalLight normal2 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[1][13]), .nBottom(GrnPixels[3][13]), .lightOn(GrnPixels[2][13]));
	normalLight normal3 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[2][13]), .nBottom(GrnPixels[4][13]), .lightOn(GrnPixels[3][13]));
	normalLight normal4 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[3][13]), .nBottom(GrnPixels[5][13]), .lightOn(GrnPixels[4][13]));
	normalLight normal5 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[4][13]), .nBottom(GrnPixels[6][13]), .lightOn(GrnPixels[5][13]));
	normalLight normal6 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[5][13]), .nBottom(GrnPixels[7][13]), .lightOn(GrnPixels[6][13]));//6
	
	centerLight center7 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[6][13]), .nBottom(GrnPixels[8][13]), .lightOn(GrnPixels[7][13]));//7
	
	normalLight normal8 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[7][13]), .nBottom(GrnPixels[9][13]), .lightOn(GrnPixels[8][13]));//8
	normalLight normal9 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[8][13]), .nBottom(GrnPixels[10][13]), .lightOn(GrnPixels[9][13]));
	normalLight normal10 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[9][13]), .nBottom(GrnPixels[11][13]), .lightOn(GrnPixels[10][13]));
	normalLight normal11 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[10][13]), .nBottom(GrnPixels[12][13]), .lightOn(GrnPixels[11][13]));
	normalLight normal12 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[11][13]), .nBottom(GrnPixels[13][13]), .lightOn(GrnPixels[12][13]));
	normalLight normal13 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[12][13]), .nBottom(GrnPixels[14][13]), .lightOn(GrnPixels[13][13]));
	normalLight normal14 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[13][13]), .nBottom(GrnPixels[15][13]), .lightOn(GrnPixels[14][13]));
	normalLight normal15 (.Clock(birdSelect), .Reset(reset| death| outofbounddeath), .up(stablePressed), .bottom(constantDown), .nUp(GrnPixels[14][13]), .nBottom(1'b0), .lightOn(GrnPixels[15][13]));//15
	

	
	// These modules are dealing with the win conditions and the 9-9-9 score counter
	winCondition(.Clock(clkSelect), .Reset(reset| death | outofbounddeath), .bird(GrnPixels), .pipes(RedPixels), .failed(death));// when green(bird) colide with red(pipes), gameover
	countScore score (.Clock(clkSelect), .Reset(reset| death | outofbounddeath), .death, .outofbounddeath, .hundredsDigit(hundreds), .tensDigit(tens), .unitsDigit(units));// Score up to 999
	Sevensegment Hex0 (.number(units), .Hex(HEX0));
	Sevensegment Hex1 (.number(tens), .Hex(HEX1));
	Sevensegment Hex2 (.number(hundreds), .Hex(HEX2));

	assign HEX3 =7'b1111111;//1 is off, 0 is on
	assign HEX4 =7'b1111111;
	assign HEX5 =7'b1111111;
	

	
endmodule


module DE1_SoC_testbench();
	
	// Testbench inputs and outputs.
	logic CLOCK_50;
	logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
	logic [9:0] LEDR;
	logic [3:0] KEY;
	logic [9:0] SW;
	logic [35:0] GPIO_1;
	
	// Instantiate the DE1_SoC module
	DE1_SoC dut(.CLOCK_50, .HEX0, .HEX1, .HEX2, .HEX3, .HEX4, .HEX5, .KEY, .LEDR, .SW, .GPIO_1);
	
	// Set up clock
	parameter CLOCK_PERIOD = 100;
	initial begin
		CLOCK_50 <= 0;
		forever #(CLOCK_PERIOD/2) CLOCK_50 <= ~CLOCK_50;
	end
	
	// Generates two possibilities: player1 wins and player2 wins.
	initial begin
	
		SW[9] <= 1;											@(posedge CLOCK_50);
		SW[9] <= 0;											@(posedge CLOCK_50);
		
		
						
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
																@(posedge CLOCK_50);
											   repeat(30) @(posedge CLOCK_50);
																
		

																
		$stop;
	end
endmodule

